PK   f�V{� l>  @    cirkitFile.json͝[s�ؕ��J�y]g���3�U��IWe*�`�X�H�Y#���˸���lP�)B�o%�T'�	,~\<X�q��4�-]�.��������n�����b�~�[��<��t1���]췋_vˏ�G�?����?>�Ǘ��ru���,���dvm��2W��Ɨ�"���zRM�����z�i��ͻ��+XX!-,+|��j����v}�_L�鼾����$���z5�L��qyyu]�E��,˼��{���ލw��M��^|��,w��y�Q�
[QD�(bV߬�]���[Q�GfT!-�0CT!-�0CT!-&a��BZL�Q�����
i1�DDyG�Z����d|�Z��U1������x�����u�w6[X̄y�L?]�%2E�UG��"z����,��H>����Oa�L?E�%2E�$����DX"S�Oa�L\�K���xf�%2E4�,.�)������Kd�xv�%2E<;��"��a�L�ΰD��ggX"Sĳ3,�k�xv�%2E<;��"��a�Lܖ�gg�ΰD��ggX"Sĳ3,�)������Kd�xv�%Ң�ggX"Sĳ3,�)������Kd
�n<;�xv�%2E<;��"��a�L�ΰD��ggX"-�xv�%2E<;��"��a�L�ΰD��ggX"S ?�ų��ggX"Sĳ3,�)������K��$��a�L�ΰD��ggKb����3�������/�!�"@R�H��	&w�`1���{��EL��Y��ar��I�z�(�E�1�~6k��U%�|ɎZ��X�\5��U�w(��t�����f�C錥��7�w�;��X�����MY�P:c��b�z7c�C錥K�9�ݜ��3�Ο�d�3�n0��`>r���M���N.O��7��`>j��2X>���y_�?��`���'�a��j��3�ϟ����+��`>:��:X>����v�?��`���'�a����3����������3��gA�����g0��߀�����`>�y��,��|>g��?X>��|��\�|��<%�?��`���V�p�����s�`�����3��g������g0��ǃҀ���`>�I��,��|>��?X>��|�&�����\�p�Q���g0�Ϙ������`>����,��|>K��?X>��|~5�\�|���p�?��`���9�\�|��l|�?��`���>�p�����`�����3��{7���3=�p�Q��G�,��|�/��?X>�����\�|�y��?��`����*�p�����}aX�j��`���6�p�����x`�����3�ϻ�����g0��?������`>���G�6�����G�5\�|�y�,�?��`���>_�p������`�����3��{���M����3�ϻ������g0�����������lYw��p��W��O���wܻl�7}�����b�t�ȁ$��O�~ڵt���F�~�'t�`����/4��5�"o_�~z��!�Z,m�����Z�l�����Zlhk!�����ů�������E��������˃㯵���@�y�~+^��p�1M�p�z����͟9h�-��:��y�g��>�?s������������<�[������M������X췋���v7z�)2���?���匇�w��<ղЏ?Ɖ�"*\�f��Pň
����5H(y�2D�P�f� ����AB�O$���AB~������u*bDs,!�Ц���WZWWK2a�mP��tX�b²۰�Rskb��۰ ��Rs	b�2ܰ��Rs�b�r��r�RJ�-9�����r�RJͭC�	���qJ)5�8!&,�,�)��܊���/���Rs�b�r��r�RJͭm�	���qJ��`LX��X�SJޠc�r��r�R�F��%�㔒7|��������1Ƅ�x��8���1&�8wS��
�qJ�'OcLX�WX�SJ>�c�r��r�R�ɨ�O?X��X�SJ>ic�r��r�R��}��&��&��5�㔒O������|Ƅ���qJ�'�`LX�O��R
O�x��'�>9��w��`%|=�W��z:��q��
����η�U��`�'X	N�@��xU���5�]_O�D0(XM��$��v�`P���5_�H|=�*�8�`5	kZ����UA_�&aM����*諂�$�iqڗW}U���՟	�k�*�4����g�5ފ�.Q٥��LSx���1�ih�Ys����KBkZf^㭦�К�֟��x���$����9o5����4�>C㭦�К���h��TdZ��������LBkZ���aAS�IhMC�s�4�j�2	�ih}Ε�[M]&�5���x���$����9po5u���4�>�O㭦.�К���$j���eZ����J����LBkZ�#��VS�IhMC�s]5�j�2	�ih}ή��$M]&�5��=�x���$����9�o5u���4�>\��iE�㊚����e��.�К����k���eZ��z�����LBkZ�VS�IhMC�=4�j�2	�ih�w��[M]&�5����x[i�2	�ih����[M]&�5��D�x���$�����.o5u���4�ޣF�h&�h*��.�4uY���$�����Ao5u���4���H㭦.�К��{8i���eZ��z/*����LBkZ�%���eZ��zo0����LBkZ�q��VS�IhMC��4�j�2	�ih���[M]&�5����x+��!j��jM]Vk�2	�ih����[M]&�5��d�x���$����ޒo5u���4��#S��DS�IhMC�>5�j�2	�ih�g��[M]&��~�״��t;P��7�@��n�U�>��.�U::oTize�{xT��n=P���@���U:z>u��eF�â��%m��4㷽��Pf w��:T��]k��aq�ʞCS��]�g�aB�k�ʡ2�(�Zr�3��V\*Ì�u��u�Qܵz��L5��W�b����quU�Ɨ�r>./��˲���e�㪦������R���r���G����G�>{��r�`�r�X�r�P�r�H�5���I]K��9>�%s<�?7:��vq�_�ףן��_�]�]��w˛c��b@B���JM�!D�Pjb!��R�$���F� ��D?B	��4�AB�9%!D�PjNo$��J&"���b�mÂ�RJ�+�	�n�RJ�;0�߆8����&,�qJ)�Z1LX�X�SJ�p?�a⮿�p,�,�)�t�m�0a9^`9N)��M�	���qJ)n�2LX�X�SJ�p�)Ǳ/����}���I�n�`9^b9N)y��	���qJ�۪`LX��X�SJ��c�r��r�R����㔒�)���{��Mq,�+,�)%�N�1a9^a9N)��e�	��
�qJɧ�b?�`9^c9N)��L�	���qJɧbLܯ��ϛX��X�SJ>mc�r��r�R�iB��,�)%���1a9>�r�Ki���&Z�0P5	�IXӢ5}�V}U���5-ZS�hU�W�IXӢ�N�V}U���5�]_[�$�&a��A_[]$�&a��(_[$�&aM�V�Z�U�jִh���UA_�&aM�V�Z�U�jV&XSh*.	�ih��f����KTvi�.�^���$����g�5�j�/	�ih��y���
LBkZ�_㭦
�К���0h��TbZ���\���jLBkZ�S��VS�IhMC�sc4�j�2	�ih}���M]&�5��U�x���$����9WoE���~��e��.+4u���4�>N㭦.�К����i���eZ����D����LBkZ�[��VS�IhMC�sD5�j�2	�ih}���[M]&�5����<����$������o5u���4�>�Z㭦.�К���k�=�(z\QS�������eZ����|����LBkZ�1��VS�IhMC�4�j�2	�ih���[M]&�5����x���$����o+M]&�5���x���$�����(o5u���4���E㭦.�К��{�h��$M%��e��.�4u���4��3H㭦.�К��{i���eZ��z'����LBkZ�E��VS�IhMC�=�$�֚�LBkZ���VS�IhMC�=�4�j�2	�ih�W��[M]&�5����x���$�����yoE]>Dm>4uY���jM]&�5��2�x���$������o5u���4��[R㭦.�К��{dJ��h�2	�ih�ק�[M]&�5��,�x���$�֏v�R��n�t�����Mv�JG�*���t������z�JG?�*��t�|:��ˌޮE_��0�kiա2��Z�t�3���	*Ì��8��@̌�U*��0��k-ȡ2�(�Zqq�3���5z�eFq��G2�t^_͊��r���U�_�������.ˢ^N�e���>*������㩏��é�������������c����C����#�ר�/3z{\���a�������_\mo���f���uu1�m�[�->�,�֫��v�ݭֻ��7o���fû���T�W���B�/��H^����7�@�	�(bNQ'��E���	*6&,��e����i�0�y��}��K������_ޮ���7��	�w����~h.����9��sN=O0���@q_�'"��|�8-�!�g'f�FORE�\�g��~�����n�ܯs}�������b�]�oV�ן"�^."_��%RsO$=�'t�[��*�P�an�b��_a����	R�%Rs�(H�H�� EX"5w��a����
R�%Rs�����$�Q�F��q�t��w�N�����h�F:�R�r 	k@��5���(���l\#~,�r Ik@��5����(��q�t��<�A\�y�H���@�@��5�ᡁ(����q�txl!��i�i\#��r yZy�H�G7�@��@��5��'��i	�i\��C@��@��5�� ��i	�i\���@�V@��5�O��i�i\��o�U�*����q�p yZy���: ����q������4��@  Ok O��c� ~�"~���4���� Ok O�>� �t�i\��%@�N�<mk��/k�t|L�5g�D>E�Mr�ڸAw[�՟{%$�Z��C�lMP�����g7Ƶ6n��z�qz�pd��˵
�_�X��|��kؿV����e�������^����̗��]���g0_Z��sqz�,��|i�����!��|��#����^�Mh4�?�I{�%xUB�%F�%�^�Mh4�?K{HW#0�ф�L/�!]���F��ȴ�tUM��R�ҕ	Lh4�?N{HW'0�ф�;�!]���F�����t�M�s���t�M��h�:&4���l��u
Lh4��7�=����hB�+C{H�)0�ф>χ���S`B�	}��!]���F��*�C�N�	�&��a��t�M���h�:&4�������u
Lh4��'�=����hB�I{H�)0�ф>�������SJ�N)�:&4������u
Lh4����=����hB��L{H�)0�ф>����S`B�	}�8�!]���F�\w�Ê�S`B�	}�>�!]���Fz��C�N�	�&����t�M�h�(�T�N��:�����hB�A{H�)0�ф�����S`B�	��	�!]���Fz�C�N�	�&�2��5]���Fz��C�N�	�&��=��t�M�}�h�:&4��{&��u
Lh4��{�=�g�����:��딚�S`B�	���!]���Fz�0�C�N�	�&��f��t�M��`'t�M�}�h�:&4��{���u
Lh�.���8tq����~����}�����c8u'�Z�M���J:p�V7с����]����Ē�UD�[G��#���P�� m�=6T :L۫}M��8m��5T ����
DGb{��ё�^�i�@t$��Iz>�����D��~��b�����F��=Z�*�;���=w��[i��٩��sP���;~������g�玞^c/<x�GO{�ء��x/�Ø�|1���f�K�g�;_۽O��^����_����ǜ�L?X&��i�w������з4��|[�ͷ6��|{���(|����=
ߣ�=
ߣ�=
ߣ�=
ߣ�=r���o�� �]v��`��z�-�j~�V}�����F��=��ц�\�v��|�x���bCg��g�s��~��)3�يs���~o�/.TlO|�:�i桫�P%zQ�������r}�IՎ�����kD�_*^*�/�/�헪����K��K����77�#�7������n��F/�'y�/�kw�^ث��?UY,�W��y��Y_����W���o��ߗ�e~�O�_���~\���usV�����ǇB��n�����=�]~�?���_�7�����L�Dv��������o���e�������:�x���cs���Y�����7��j�z�?G�">,oﯗW���z���fG$����v�d����f�}x3.��մ>��Ŭ(^��N'�)V�u����xZ�|���r<�,��L�iU��͗=����a�^?��n����ft�1���fwu�~�3`]������|��|����g>����i�+6��Ǧ��L:��:���WR�ڬk�i�u�U�e�d'���4��?L�_��RMӯ��v�>_^�I�+�k�u�c��}����Wʖ_^i7_^i7��������������w�/�k�������_m��X��Ǉ���ɩ͵r2I�C���׻���O?ݮ�}��I������&�W�bfE����8�&�y=Ou1.g+O��j<���㺬�����zZ��Oqto�y�p���E�l��)5'��z8־�T������I��i�����R��e��ᵣ7���n����f�"͎ �|��/�_ޠ�(��++뺘��޲��jb�|j�;6(�;Nf�#|ݠ,R:�`���@6�z}�jjդ�^�9�����T�7(�WŤ�M��c����/>}����]5-�W�dV~���~ݳ��]5�~�������[���z���!����Y�߻B������/�}����޿����#y���z�^�������z�����o����;����6G��v�v�����6�������m>d���ϛ۟V�K/.�����	�h��H��D�z��������^��7ڟ޾};��]��/����;���o��O.<�/_�oq��f�T��v9T����v���fգ������v�9��ǣ�����QV�FY>q�����/�CG��K��Qv�ټcTL_�٤H��Xk����@yf��vnX}���_�����GV=?�^�:tLU�.�_�`Z_�k�����9�sL�7�NK�Ƨr�$:��@��I�(y�Y߬�q���\V������x��[�z���f_*�3Y1p�C�)�;�1��A9��Hy=:�:"�d����i]]-�>�����B_��/���{]��l�p��lZ�̦�����;U�~��39�2��z:8�Gt���
��W9U�)�Q���:���s1U���N��e�i�/�o�pg�l����>qwJ�6���T��
�(fTu\ܜn6}2Z��u�A��luP~�|ss��.���fy���k������������?����c��<���PK
   f�V{� l>  @                  cirkitFile.jsonPK      =   k    