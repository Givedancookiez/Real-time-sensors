PK   w �V���i�  B    cirkitFile.json�]o"Y�E�J�~5V����53%�CO�ԣ����*�8M��1���}O�L�a"��UҔTݕI�a������i�[�����lw��ϫ��f{7���b�~�[��x�������n����->�]}�?���}\��w���z�Ι�V�z���xQ���in��Y���|]��dYOo��l���޼���
���-Ux:�f����nu��O�ɬ�����u��˛j9�ήg���f]y��E:��s���ڍw��m����.v��o���QL
K�G��cR�ORܭ~
J���(�#3Z!��a�h�l^���yf�V��0C�B6�����,b�s�x:w�-�j�X�������"�[�7����\T�r�.�:�	��'E��*\"Q�>���[0�~B�?�,j�/�(���"�.�(���"�!.�(���"�A.�(��k�iZ��p�D5>��Hq��Hq��Hq��Hq���|j��{g��p�D��p�D��p�����.�(��.�(��.�(��%��YĽ3\"QĽ3\"QĽ3\"QĽ3\"QĽ3\"QĽ3\"��q��Hq��Hq��Hq��H���q�,��.�(��.�(��.�(��.�(��.�ͫ�w�K$��w�K$��w�K$��w�K$��w�K$
�'��wVq��Hq��Hq��Hq����u�;�%E�;�%E�;[%��ؐ�����ow�~�r���=�<�bmU�r�Wʺ߳o�����6k�6��|Nҵ�*����1��6k���T�|��Z��X���X�JV;��X�4ob��X�P:c���ծf�C錥��V�	�Jg,]6���MY�P:c����n�j��K�w`����3�������	N�tbp<1to0��|~�,��2X>����_X?8i�|���ʰ~p�`���a���������������3���l�����g0�ߓ����`>_M =���`>_����`>_�����`>_{����`>_5����`>_�����`>_�����`>_c����`>_����`>_�����`>_�ߤ���`>_K����`>_	����`>_�	�G�eE�f���?X>��|�,��?X>��|�/��?X>��|�2��?X>��|�5��?X>��|m8��?X>��|U;�_	���`>_�����`>�$ ����`>� ����`>�� �G����z�����G	���`>�����`>������`>�R����`>�����`>���W����3��{�������3�ϻ�������3���������3��; ������3��{7��ѫ����p����Q����3���e������3��;}������3��{�������3�ϻ����p�`���p�~p�`���v�~p�`����������l7xsE�u��m�bO>�<�q�����ߵ��v�au��ǭQ�~��t����H�^/������[w=��a���Gn�������;�[�^�wk����t����}��:����uz�U���߰��ำ��tç4G3�Jp7 ���ݡ�����ֈC�^�����*Z[ =?��A;nm�7���!�6����f
�w���$�s����v~����FW�"�x�9k�y�����P!�7����ǉ�"ʽ�Mg����QA�kP�f�y�*�l8�A����"�P�=Cj��g��B�F��?�׫*�cD3�!1Ӧ*6�O�V��L�o䷆U:l�1a�m�yS���CL�f�T��F��ᆙ8U鰉<Ą�x��8U��<��Ϳ1�*6���0�1�*6���0�1�*6���0�1�*6���0/0�*6���0/0�*e�.�����T����b�|��|���$0&���ǩJ�� c�|��|����1&��K�ǩJ��c���|��|��䋇1&��K�ǩJ��c�|��|���1��~0�0�*��A�	��
�q��/nØ�_7��71�0�*��&�	��
�q��/���0�1�*�B�	����J�[O���'��m9���Y�
�	VB��uE��ǫ�ڬpUP���FxUp�*X�+��q�*8^�&aM�K��q�F�IX�<H��q�F�IX�E��qWF�IX��q��*����$�����^�U�j�l~ܗ�
�`5	��,�)�4����{�5ڊR�(vir�i��)ҌihMC���k�դ/	�ih��y���&�5�����V��$����5m5ILBkZ_���V��$����5%m5�LBkZ_��V��$����5>�4�LBkZ_���V��$����5Wm5�LBkZ_;��V��$����5pm5�LBkZ_˧�V��$����5�m5�LBkZ_[��V��$����5�m5�LBkZ_��V��$����5���4�LBkZ_{��V��$����5�m5�LBkZ_��Vt���vEM.+4����2	�ih}m�F[M.�К��{h���2	�ih�W�F[M.�К��{>h���2	�ih�w�F[M.�К��{pH�-5�LBkZ�%��V��$�����(m5�LBkZ���V��$����5mE+�DK�4����R��$�����Am5�LBkZ�}��V��$����Nm5�LBkZ�E��V��$�����Zm+M.�К��{�i���2	�ih�ǙF[M.�К��{�i���2	�ih��F[M.�К��{�i�u�����J��*M.�К��{j���2	�ih�'�F[M.�К��{Kj���2	�ih�G�D�Z��$����^�m5�LBkZ�Y��V��$�֏�i��I9�U7�|����qyS-����l\\߬�"����ڇy`��M�V��8y`���w{ցU::o�r����t`�����t��X�����*=���:h�vtVZ����2}臖9;�{mAV�^U�
ܫ�Y}{U9+o�*����V9k�����^U��C�*g�ߨ�/3z��[�2��=��k����0#�k�e�1ܵ���2�(�ګwhȃ���vhƆ���Z�>7��Wf�l����3�o����~5���Tw��>��V����9����BY33@��BY3�@��BY3cA��BY3�A��BY3�B��BY3+C��BY3�C��BY3[D��BY3�D��B�a�X$�ڜmc�m�qS���d�a¼�0�*e��0a�m��S��C�a�07�ĩJ�!z1L��瘏S��C(d���77�|<�|����/Ä�x��8U);�r�	���q����0�1�*y�&,�c>^`>NU�A�M
�U
����T%o�1a>^`>NU��!����T%oU�1a>^b>NU����%��T%_��1q߉s_�c>^b>NU�%���%��T%_��1a>^b>NU�%��O?��W��S�|	"Ƅ�x��8Uɗ�aLܯ��ϛ��W��S�|iƄ�x��8Uɗ�`L��ט�S�|�Ƅ�x��xW���(Z�t誇�@U����5�����UA]�&a���9tUPW�IX�y�e]�U�j֔�$���% 
(XM�A][��&aMs���.	�
V��f�V��*����$�ټ���
�`5	k6o�F����*XM���k��&qIhMC��6k��.Q���.�/�$/	�ih�^s����%�5��3��V��$����{�5�jR���4���A��&�IhMC�k14�jҘ��4���D��&�IhMC�kc4�jR���4���G�Â&�IhMC�k�4�jr���4���J���1�Ob�\�krY��eZ���8���\&�5����h��eZ����D���\&�5����h��eZ���Q���\&�5��u�h��eZ����]͍I�\&�5��=�h��eZ���j���\&�5���h+�[Qt��&��\Vhr���4��6_��&�IhMC�=4�jr���4��+A��&�IhMC�=4�jr���4�޻B��&�IhMC�=8$ږ�\&�5���h��eZ��zO���\&�5��v�h��eZ��z�����d��d�\VjrY��eZ��z� ���\&�5��>�h��eZ��z'���\&�5����h��eZ��zO-���&�IhMC��4�jr���4���L��&�IhMC��4�jr���4��sN��&�IhMC��4ڊ�|��|hrY��e�&�IhMC�5�jr���4�ޓQ��&�IhMC�%5�jr���4��#S�m��eZ��z�O���\&�5��,�h��eZ�G��W���̪�i>^]�ٸ������z6.�o�E�W�zQt��<�JGoځU:������{`�����t��X�����*��V�� =�JG�硣������uhf�vm�:p+��
��rV�~��#U��۫
��Y{�U�=��r�zU9k�����~����=o��0����͒��a�pז�C�0��k�ߡ�ǌ��u��aFq�&�C�0��k�ءe�Q�bC���?��o����|��utU^�~��V�󏷋��r���ow��nt�����e׶^���r�JO:)ǳ��f�X����*�;��O�P�:
��.����H<yEH�	I�x���63���R ��qJ�1%�yL���u�/Z�Ƅ����=�,<"�����-<f�g/���;��Xu�I��!�!��CW3$��޽��[}���>�w�S�o��s��Ä��!� �qh.����!��kf#'~�II\�������uf*q������yB�����ã��q|5D6��~��r��w��D�i��[zO�����3��|����~�دFW_��]������a�]}���W�����Kdͯc��BS���mA���=�|�*��W�D�����Ț���Y��c�"\"k~�R�Kd�o�A�p�������M���F-p�x���[�:e0[{�5�Ï�Q�a��x����v�pYl6^#;��� �� ����?�G9 {�{���7D9��+����6�(�9����F�(�9����V�(�9���j� �� �4^�[X�����kxkd�����xo�p ~Z ~��\�O�O�5�E(��i	�i����8 ?-?��� �*�*�%���V� ���4^�ە������kx,���O+�O�5����i�i����8�ߨ�� ?� ?����) ���ޒ� ���4^�[= ��ր��k�o�i�t����|)om������j ��M(�� ��q�z����\���3t��������V�E�2Y>��RV��k�V�^��`�47��k�O�^��`�4���k�H�^��`�l�j���C�c���歖�\=D?��`�l�jk��C�c���[a���Mh4�߮Ik��<�б��\b�L�hB�	��XZC:���F�=���t"�	�&���i�TM��R���&4����5��	Lh4���NkH'��hB���֐N)0�ф�v��ޚ�)0�ф��֐�)0�ф�f�֐�)0�ф�ބ֐�)0�ф�V�֐�)0�ф�·֐�)0�ф�F�֐�)0�ф���֐�)0�ф�6�֐�)0�ф���֐�)0�ф�&��!��)0�ф���֐�)0�ф��֐�)0�ф����������)�S
:���F��YZC:���F��_ZC:���F��eZC:���F��kZC:���F�zqZC:���F�ZwXÒ�)0�ф�N�֐�)0�ф�c�֐�)0�ф��֐�)0�ф�ہ�_��/E�sJI甒�)0�ф�S�֐�)0�ф��֐�)0�ф�˄֐�)0�фއ�֐�)0�ф�Cְ�s
Lh4����5�s
Lh4���5�s
Lh4���5�s
Lh4��L�5�s
Lh4��{�5�W�����R�9��s
Lh4��٢5�s
Lh4���5�s
Lh4��7�5�s
Lh4��f�5��M�}�h�M�=�h��9;��#�v��u�wk~������_�vm`�V���{.�����r�ާ�o�,x~�����[=B�����mu�Z��Nsh�V_�^��vw}E�~���E�^�"`����!<�������\Ľ��"�u�+q����h'>t�H��l��ך����]
�������CD�i{'���N����uCDͲ�M�������n�~bJ��b�Tg��m������}>�GWoFn ~��d�g�>�s�:�;I�Nӿ�)�5��懚���w����3����7?���3r?#oj����������A}R�� ��j��Vz�Xp�¾�{��P(<����V_[,2�^�Q�l��2��E޸��~5U���Bi4d|���x1ç=����8�+1��}2������vq��u�j���?W�?�6�k�y�h?T>>T����e�e���!������@�ܭ��������F�Lb�_����.g���X5��/y'���z�o���_G���/���l����q�����7��3���;�?I���ns�S��n����^�~^�>����v}�6�}����������[*:�Z/n�W��������������V���٭���}z�]���{X/n����g~��_����a���w�?'��8U�J�{��l� oƕUe=���S˫� n�Tu��I�z:�fY�����f�Ȗ��Z/�UQ�̖���z�c8�u�����9�f<�mzMw�ŁeԼ�����nnW�o�q9�\V	����?dY3��<����i�<T�/�gM��,��U�YV�{�dey8mR>���9>Ϧ� ��.mbY��	��bV\ZQU��zz�ʲ��f���:��3������aE�e��]V	�&]�O/'V���*��I��uy��8f�y]M'y�q@�����?{��/Ǖ��p@vY��⩀?�y�g����a���c��?��I�K7���Y6����g>�]�&u�ި�;[]L�/˞����Z�f�z}3����U�X��:�^/g��E==�X{�����c�R5�8��tq1�6����K�T��#Ծ>�g����`��@~8%�ۏ���G��if��R���R8<P~}�nN�N��S��)���Ϛ3ʯ��W�S�ɣY�_țS�����pFѮUN��֤9%�L�|}dڜ�^��ev8%�����^|��i�Ӈ�^���Nx���;p���;x���8}\k�>�=O��';q�>�}!��;�>�>�-�o?�s~��t�6��W�q������Y��{�l����W������ٗ觞�=>����ː�������w����lV��w��{�~z�>	n�������?����vt�69�b��qs�òy($�z���jC�hJ����,����z����w�����~�n��?.��Z�޾};�����?�o>���o����~1���_fY�����a�$pX��0�69sػ�oG�� ��K� ���^<zt0����au~|��ߦ��|W�o�yE�{�s�+�oz{g!�L��/��W<��:-�}�dLE�wU�1�RN�G�\��Vgǃ��۟�ʛ�џ(���~���������9S9:����n1�0����J�?ި����tX��o�����8:�Ο��O��g�����z���03΅
�p��&T|�`��3���=~�|�]��Uu�	��Í���S*lA52��,��auqz"��{�އ�����?���l�4��X���	��S���'��i��6/m��a���a�M������_5�z|�m��Q���ټ�i�{��<lj�~�e=ktz�u|Q�_zono����b��m��x&�����[-���{X�~����~���_��ϣ��PK
   w �V���i�  B                  cirkitFile.jsonPK      =   �    